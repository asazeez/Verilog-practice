library verilog;
use verilog.vl_types.all;
entity lab1block_vlg_vec_tst is
end lab1block_vlg_vec_tst;
