library verilog;
use verilog.vl_types.all;
entity asu_vlg_vec_tst is
end asu_vlg_vec_tst;
