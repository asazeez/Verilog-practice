library verilog;
use verilog.vl_types.all;
entity orgate_vlg_vec_tst is
end orgate_vlg_vec_tst;
