library verilog;
use verilog.vl_types.all;
entity fullasublock_vlg_vec_tst is
end fullasublock_vlg_vec_tst;
