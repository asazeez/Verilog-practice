library verilog;
use verilog.vl_types.all;
entity orgate_vlg_check_tst is
    port(
        pin_name3       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end orgate_vlg_check_tst;
